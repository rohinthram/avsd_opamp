
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

* Stage 1 - Differential amplifier
xm1 net-_m1-pad1_ in1 net-_m1-pad3_ net-_m1-pad3_ sky130_fd_pr__nfet_01v8 l=1 w=1.79
xm2 out1 in2 net-_m1-pad3_ net-_m1-pad3_ sky130_fd_pr__nfet_01v8 l=1 w=1.79
xm3 net-_m1-pad1_ net-_m1-pad1_ vdd vdd sky130_fd_pr__pfet_01v8 l=1 w=10
xm4 out1 net-_m1-pad1_ vdd vdd sky130_fd_pr__pfet_01v8 l=1 w=10

* Current Mirror
xm5 net-_m1-pad3_ ref vss vss sky130_fd_pr__nfet_01v8 l=1 w=20
xm6 ref ref vss vss sky130_fd_pr__nfet_01v8 l=1 w=10

* Stage 2 - PMOS Common Source Amplifier
xm7 out2 out1 vdd vdd sky130_fd_pr__pfet_01v8 l=1 w=62.83
xm8 out2 ref vss vss sky130_fd_pr__nfet_01v8 l=1 w=62.83


* Circuit Bias
v1  vdd gnd dc 1
v2  vss gnd dc -1
xR1 vdd ref gnd sky130_fd_pr__res_high_po_0p69 l=100


v3 in1 gnd ac 1
v4 in2 gnd ac 1

*Simulation Command
*.tran 0.1e-3 10e-3 0
.ac dec 101 1 1g

* ngspice control statements
.control

run
print allv > plot_data_v.txt
print alli > plot_data_i.txt

*For Transient Analysis
*plot v(in1)
*plot v(in2)
*plot v(out2)

*For AC Analysis
plot db(V(out2)/V(in1))

let gain = db(V(out2)/V(in1))
let max_gain = maximum(gain)

print max_gain

.endc
*results
*Acm = -8.399db

.end
