* SPICE3 file created from avsd_opamp_layout.ext - technology: sky130A

.option scale=10000u

X0 a_181_n17# in1 a_n28_306# vss sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=179 l=100
X1 vss a_n675_n1020# out2 vss sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=6289 l=100
X2 vss a_n675_n1020# a_n675_n1020# vss sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1001 l=100
X3 out2 a_582_n17# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=6289 l=100
X4 a_n1220_n998# a_n1049_1511# vss sky130_fd_pr__res_generic_nd w=27 l=2492
X5 a_582_n17# a_n28_306# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1001 l=100
X6 a_n1220_n998# vdd vss sky130_fd_pr__res_generic_nd w=27 l=2492
X7 a_n883_n1009# a_n1049_1511# vss sky130_fd_pr__res_generic_nd w=27 l=2492
X8 vdd a_n28_306# a_n28_306# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1001 l=100
X9 a_582_n17# in2 a_181_n17# vss sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=179 l=100
X10 a_n675_n1020# a_n883_n1009# vss sky130_fd_pr__res_generic_nd w=26 l=2494
X11 vss a_n675_n1020# a_181_n17# vss sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2002 l=100
C0 vss vss 5.09fF
C1 a_n675_n1020# vss 5.61fF
C2 a_n883_n1009# vss 3.88fF
C3 vdd vss 125.23fF
