magic
tech sky130A
timestamp 1629189414
<< nwell >>
rect -107 244 1438 6840
<< nmos >>
rect 81 -17 181 162
rect 482 -17 582 162
rect -187 -2092 -87 -1091
rect 347 -2232 447 -230
rect 1643 -2149 1743 4140
<< pmos >>
rect 77 306 177 1307
rect 506 306 606 1307
rect 936 425 1036 6714
<< ndiff >>
rect 1537 3857 1643 4140
rect 1538 2118 1643 3857
rect 1538 2078 1563 2118
rect 1604 2078 1643 2118
rect 1538 2029 1643 2078
rect 1538 1989 1563 2029
rect 1604 1989 1643 2029
rect -21 138 81 162
rect -21 98 1 138
rect 42 98 81 138
rect -21 49 81 98
rect -21 9 1 49
rect 42 9 81 49
rect -21 -17 81 9
rect 181 138 291 162
rect 181 98 220 138
rect 261 98 291 138
rect 181 43 291 98
rect 181 3 216 43
rect 257 3 291 43
rect 181 -17 291 3
rect 380 138 482 162
rect 380 98 402 138
rect 443 98 482 138
rect 380 49 482 98
rect 380 9 402 49
rect 443 9 482 49
rect 380 -17 482 9
rect 582 138 692 162
rect 582 98 621 138
rect 662 98 692 138
rect 582 43 692 98
rect 582 3 617 43
rect 658 3 692 43
rect 582 -17 692 3
rect 1538 116 1643 1989
rect 1538 76 1563 116
rect 1604 76 1643 116
rect 1538 27 1643 76
rect 1538 -13 1563 27
rect 1604 -13 1643 27
rect 242 -309 347 -230
rect 242 -349 278 -309
rect 319 -349 347 -309
rect -292 -1153 -187 -1091
rect -292 -1193 -255 -1153
rect -214 -1193 -187 -1153
rect -292 -1829 -187 -1193
rect -292 -1869 -267 -1829
rect -226 -1869 -187 -1829
rect -292 -1918 -187 -1869
rect -292 -1958 -267 -1918
rect -226 -1958 -187 -1918
rect -292 -2092 -187 -1958
rect -87 -1829 26 -1091
rect -87 -1869 -48 -1829
rect -7 -1869 26 -1829
rect -87 -1924 26 -1869
rect -87 -1964 -52 -1924
rect -11 -1964 26 -1924
rect -87 -2092 26 -1964
rect 242 -1969 347 -349
rect 242 -2009 267 -1969
rect 308 -2009 347 -1969
rect 242 -2058 347 -2009
rect 242 -2098 267 -2058
rect 308 -2098 347 -2058
rect 242 -2232 347 -2098
rect 447 -1969 560 -230
rect 447 -2009 486 -1969
rect 527 -2009 560 -1969
rect 447 -2064 560 -2009
rect 447 -2104 482 -2064
rect 523 -2104 560 -2064
rect 447 -2232 560 -2104
rect 1538 -1886 1643 -13
rect 1538 -1926 1563 -1886
rect 1604 -1926 1643 -1886
rect 1538 -1975 1643 -1926
rect 1538 -2015 1563 -1975
rect 1604 -2015 1643 -1975
rect 1538 -2149 1643 -2015
rect 1743 2118 1856 4140
rect 1743 2078 1782 2118
rect 1823 2078 1856 2118
rect 1743 2023 1856 2078
rect 1743 1983 1778 2023
rect 1819 1983 1856 2023
rect 1743 116 1856 1983
rect 1743 76 1782 116
rect 1823 76 1856 116
rect 1743 21 1856 76
rect 1743 -19 1778 21
rect 1819 -19 1856 21
rect 1743 -1886 1856 -19
rect 1743 -1926 1782 -1886
rect 1823 -1926 1856 -1886
rect 1743 -1981 1856 -1926
rect 1743 -2021 1778 -1981
rect 1819 -2021 1856 -1981
rect 1743 -2149 1856 -2021
<< pdiff >>
rect 830 6431 936 6714
rect 831 4692 936 6431
rect 831 4652 856 4692
rect 897 4652 936 4692
rect 831 4603 936 4652
rect 831 4563 856 4603
rect 897 4563 936 4603
rect 831 2690 936 4563
rect 831 2650 856 2690
rect 897 2650 936 2690
rect 831 2601 936 2650
rect 831 2561 856 2601
rect 897 2561 936 2601
rect 831 1574 936 2561
rect 831 1534 865 1574
rect 906 1534 936 1574
rect -28 1253 77 1307
rect -28 1213 5 1253
rect 46 1213 77 1253
rect -28 569 77 1213
rect -28 529 -3 569
rect 38 529 77 569
rect -28 480 77 529
rect -28 440 -3 480
rect 38 440 77 480
rect -28 306 77 440
rect 177 1242 290 1307
rect 177 1202 215 1242
rect 256 1202 290 1242
rect 177 569 290 1202
rect 177 529 216 569
rect 257 529 290 569
rect 177 474 290 529
rect 177 434 212 474
rect 253 434 290 474
rect 177 306 290 434
rect 401 1242 506 1307
rect 401 1202 437 1242
rect 478 1202 506 1242
rect 401 569 506 1202
rect 401 529 426 569
rect 467 529 506 569
rect 401 480 506 529
rect 401 440 426 480
rect 467 440 506 480
rect 401 306 506 440
rect 606 569 719 1307
rect 606 529 645 569
rect 686 529 719 569
rect 606 474 719 529
rect 606 434 641 474
rect 682 434 719 474
rect 606 306 719 434
rect 831 688 936 1534
rect 831 648 856 688
rect 897 648 936 688
rect 831 599 936 648
rect 831 559 856 599
rect 897 559 936 599
rect 831 425 936 559
rect 1036 4692 1149 6714
rect 1036 4652 1075 4692
rect 1116 4652 1149 4692
rect 1036 4597 1149 4652
rect 1036 4557 1071 4597
rect 1112 4557 1149 4597
rect 1036 2690 1149 4557
rect 1036 2650 1075 2690
rect 1116 2650 1149 2690
rect 1036 2595 1149 2650
rect 1036 2555 1071 2595
rect 1112 2555 1149 2595
rect 1036 2109 1149 2555
rect 1036 2069 1075 2109
rect 1116 2069 1149 2109
rect 1036 688 1149 2069
rect 1036 648 1075 688
rect 1116 648 1149 688
rect 1036 593 1149 648
rect 1036 553 1071 593
rect 1112 553 1149 593
rect 1036 425 1149 553
<< ndiffc >>
rect -516 1525 -489 1556
rect -440 1511 -413 1542
rect -516 -998 -489 -967
rect -368 1514 -341 1545
rect -247 1505 -220 1536
rect -440 -1012 -413 -981
rect -368 -1009 -341 -978
rect 1563 2078 1604 2118
rect 1563 1989 1604 2029
rect 1 98 42 138
rect 1 9 42 49
rect 220 98 261 138
rect 216 3 257 43
rect 402 98 443 138
rect 402 9 443 49
rect 621 98 662 138
rect 617 3 658 43
rect 1563 76 1604 116
rect 1563 -13 1604 27
rect 278 -349 319 -309
rect -248 -1020 -221 -989
rect -255 -1193 -214 -1153
rect -267 -1869 -226 -1829
rect -267 -1958 -226 -1918
rect -48 -1869 -7 -1829
rect -52 -1964 -11 -1924
rect 267 -2009 308 -1969
rect 267 -2098 308 -2058
rect 486 -2009 527 -1969
rect 482 -2104 523 -2064
rect 1563 -1926 1604 -1886
rect 1563 -2015 1604 -1975
rect 1782 2078 1823 2118
rect 1778 1983 1819 2023
rect 1782 76 1823 116
rect 1778 -19 1819 21
rect 1782 -1926 1823 -1886
rect 1778 -2021 1819 -1981
<< pdiffc >>
rect 856 4652 897 4692
rect 856 4563 897 4603
rect 856 2650 897 2690
rect 856 2561 897 2601
rect 865 1534 906 1574
rect 5 1213 46 1253
rect -3 529 38 569
rect -3 440 38 480
rect 215 1202 256 1242
rect 216 529 257 569
rect 212 434 253 474
rect 437 1202 478 1242
rect 426 529 467 569
rect 426 440 467 480
rect 645 529 686 569
rect 641 434 682 474
rect 856 648 897 688
rect 856 559 897 599
rect 1075 4652 1116 4692
rect 1071 4557 1112 4597
rect 1075 2650 1116 2690
rect 1071 2555 1112 2595
rect 1075 2069 1116 2109
rect 1075 648 1116 688
rect 1071 553 1112 593
<< psubdiff >>
rect -184 -127 -66 -98
rect -184 -197 -169 -127
rect -99 -197 -66 -127
rect -184 -217 -66 -197
<< nsubdiff >>
rect 556 1693 594 1698
rect 527 1684 652 1693
rect 527 1654 563 1684
rect 586 1654 652 1684
rect 527 1641 652 1654
<< psubdiffcont >>
rect -169 -197 -99 -127
<< nsubdiffcont >>
rect 563 1654 586 1684
<< poly >>
rect 936 6714 1036 6737
rect 75 1422 188 1439
rect 75 1339 96 1422
rect 161 1339 188 1422
rect 75 1316 188 1339
rect 506 1421 606 1436
rect 506 1338 529 1421
rect 594 1338 606 1421
rect 77 1307 177 1316
rect 506 1307 606 1338
rect 1643 4140 1743 4163
rect 936 366 1036 425
rect 936 329 954 366
rect 986 329 1036 366
rect 936 312 1036 329
rect 77 260 177 306
rect 506 260 606 306
rect 81 162 181 196
rect 482 162 582 196
rect 81 -76 181 -17
rect 482 -25 582 -17
rect 81 -114 99 -76
rect 146 -114 181 -76
rect 81 -138 181 -114
rect 481 -70 582 -25
rect 481 -108 512 -70
rect 559 -108 582 -70
rect 481 -137 582 -108
rect 81 -139 180 -138
rect 347 -230 447 -205
rect -187 -1091 -87 -1043
rect -187 -2107 -87 -2092
rect -188 -2290 -85 -2107
rect 1643 -2162 1743 -2149
rect -188 -2325 -161 -2290
rect -107 -2325 -85 -2290
rect -188 -2370 -85 -2325
rect 347 -2283 447 -2232
rect 347 -2318 367 -2283
rect 421 -2318 447 -2283
rect 1641 -2268 1743 -2162
rect 1641 -2301 1671 -2268
rect 1719 -2301 1743 -2268
rect 1641 -2304 1743 -2301
rect 1647 -2316 1741 -2304
rect 347 -2339 447 -2318
<< polycont >>
rect 96 1339 161 1422
rect 529 1338 594 1421
rect 954 329 986 366
rect 99 -114 146 -76
rect 512 -108 559 -70
rect -161 -2325 -107 -2290
rect 367 -2318 421 -2283
rect 1671 -2301 1719 -2268
<< ndiffres >>
rect -521 1556 -484 1573
rect -521 1525 -516 1556
rect -489 1525 -484 1556
rect -521 -611 -484 1525
rect -445 1542 -408 1559
rect -445 1511 -440 1542
rect -413 1511 -408 1542
rect -521 -967 -485 -611
rect -521 -998 -516 -967
rect -489 -998 -485 -967
rect -521 -1004 -485 -998
rect -445 -625 -408 1511
rect -373 1545 -336 1562
rect -373 1514 -368 1545
rect -341 1514 -336 1545
rect -373 -622 -336 1514
rect -252 1536 -215 1553
rect -252 1505 -247 1536
rect -220 1505 -215 1536
rect -445 -981 -409 -625
rect -445 -1012 -440 -981
rect -413 -1012 -409 -981
rect -445 -1018 -409 -1012
rect -373 -978 -337 -622
rect -373 -1009 -368 -978
rect -341 -1009 -337 -978
rect -373 -1015 -337 -1009
rect -252 -631 -215 1505
rect -252 -989 -216 -631
rect -252 -1020 -248 -989
rect -221 -1020 -216 -989
rect -252 -1026 -216 -1020
<< locali >>
rect 841 4692 907 4705
rect 841 4652 856 4692
rect 897 4652 907 4692
rect 841 4634 907 4652
rect 1061 4692 1127 4705
rect 1061 4652 1075 4692
rect 1116 4652 1127 4692
rect 1061 4634 1127 4652
rect 841 4603 907 4616
rect 841 4563 856 4603
rect 897 4563 907 4603
rect 841 4545 907 4563
rect 1061 4597 1127 4617
rect 1061 4557 1071 4597
rect 1112 4557 1127 4597
rect 1061 4546 1127 4557
rect 841 2690 907 2703
rect 841 2650 856 2690
rect 897 2650 907 2690
rect 841 2632 907 2650
rect 1061 2690 1127 2703
rect 1061 2650 1075 2690
rect 1116 2650 1127 2690
rect 1061 2632 1127 2650
rect 841 2601 907 2614
rect 841 2561 856 2601
rect 897 2561 907 2601
rect 841 2543 907 2561
rect 1061 2595 1127 2615
rect 1061 2555 1071 2595
rect 1112 2555 1127 2595
rect 1061 2544 1127 2555
rect 1065 2116 1131 2129
rect 1548 2118 1614 2131
rect 1548 2116 1563 2118
rect 1065 2109 1563 2116
rect 1065 2069 1075 2109
rect 1116 2078 1563 2109
rect 1604 2078 1614 2118
rect 1116 2076 1614 2078
rect 1116 2069 1131 2076
rect 1065 2058 1131 2069
rect 1548 2060 1614 2076
rect 1768 2118 1834 2131
rect 1768 2078 1782 2118
rect 1823 2078 1834 2118
rect 1768 2060 1834 2078
rect 1548 2029 1614 2042
rect 1548 1989 1563 2029
rect 1604 1989 1614 2029
rect 1548 1971 1614 1989
rect 1768 2023 1834 2043
rect 1768 1983 1778 2023
rect 1819 1983 1834 2023
rect 1768 1972 1834 1983
rect 549 1686 681 1693
rect 549 1684 687 1686
rect 549 1680 563 1684
rect 547 1654 563 1680
rect 586 1654 687 1684
rect 547 1628 687 1654
rect -150 1617 -112 1618
rect -522 1588 -110 1617
rect -520 1561 -482 1588
rect -150 1586 -112 1588
rect -149 1564 -112 1586
rect 651 1575 687 1628
rect 850 1575 916 1587
rect 651 1574 916 1575
rect 651 1571 865 1574
rect 35 1564 865 1571
rect -371 1562 -337 1564
rect -519 1556 -484 1561
rect -519 1525 -516 1556
rect -489 1525 -484 1556
rect -519 1522 -484 1525
rect -518 1514 -484 1522
rect -443 1559 -409 1560
rect -443 1551 -408 1559
rect -371 1551 -336 1562
rect -149 1556 865 1564
rect -236 1553 -213 1555
rect -443 1545 -336 1551
rect -443 1542 -368 1545
rect -443 1511 -440 1542
rect -413 1516 -368 1542
rect -413 1511 -408 1516
rect -371 1514 -368 1516
rect -341 1514 -336 1545
rect -249 1536 -213 1553
rect -371 1511 -336 1514
rect -443 1508 -408 1511
rect -442 1500 -408 1508
rect -370 1503 -336 1511
rect -307 1533 -279 1536
rect -250 1533 -247 1536
rect -307 1505 -247 1533
rect -220 1518 -213 1536
rect -149 1552 441 1556
rect -149 1532 217 1552
rect 244 1536 441 1552
rect 468 1536 865 1556
rect 244 1534 865 1536
rect 906 1534 916 1574
rect 244 1532 916 1534
rect -149 1521 916 1532
rect -220 1505 -215 1518
rect 850 1516 916 1521
rect -307 1501 -215 1505
rect -307 852 -279 1501
rect -249 1494 -215 1501
rect 72 1438 193 1446
rect 72 1422 607 1438
rect 4 1382 41 1385
rect 72 1382 96 1422
rect 4 1349 96 1382
rect 4 1266 41 1349
rect 72 1339 96 1349
rect 161 1421 607 1422
rect 161 1339 529 1421
rect 72 1338 529 1339
rect 594 1338 607 1421
rect 72 1321 607 1338
rect 72 1315 193 1321
rect -9 1253 57 1266
rect -9 1213 5 1253
rect 46 1213 57 1253
rect -9 1195 57 1213
rect 201 1242 267 1255
rect 201 1202 215 1242
rect 256 1202 267 1242
rect 201 1184 267 1202
rect 423 1242 489 1255
rect 423 1202 437 1242
rect 478 1202 489 1242
rect 423 1184 489 1202
rect -307 836 -277 852
rect -305 474 -277 836
rect 841 688 907 701
rect 841 648 856 688
rect 897 648 907 688
rect 841 630 907 648
rect 1061 688 1127 701
rect 1061 648 1075 688
rect 1116 648 1127 688
rect 1061 630 1127 648
rect 841 599 907 612
rect -18 569 48 582
rect -18 529 -3 569
rect 38 529 48 569
rect -18 511 48 529
rect 202 569 268 582
rect 202 529 216 569
rect 257 529 268 569
rect 202 511 268 529
rect 411 569 477 582
rect 411 529 426 569
rect 467 529 477 569
rect 411 511 477 529
rect 631 569 697 582
rect 631 529 645 569
rect 686 529 697 569
rect 841 559 856 599
rect 897 559 907 599
rect 841 541 907 559
rect 1061 593 1127 613
rect 1061 553 1071 593
rect 1112 553 1127 593
rect 1061 542 1127 553
rect 631 511 697 529
rect 1071 502 1104 542
rect -309 419 -277 474
rect -18 480 48 493
rect -18 440 -3 480
rect 38 440 48 480
rect -18 422 48 440
rect 202 474 268 494
rect 202 434 212 474
rect 253 434 268 474
rect 202 423 268 434
rect 411 480 477 493
rect 411 440 426 480
rect 467 440 477 480
rect 631 474 697 494
rect 631 461 641 474
rect 411 422 477 440
rect 628 434 641 461
rect 682 434 697 474
rect 628 423 697 434
rect 1071 461 1365 502
rect 1071 428 1104 461
rect -309 -17 -278 419
rect 5 151 32 422
rect 628 217 673 423
rect 1056 372 1098 386
rect 944 366 1098 372
rect 944 329 954 366
rect 986 329 1098 366
rect 944 325 1098 329
rect 1056 237 1098 325
rect 1056 217 1080 237
rect 1170 217 1200 461
rect 628 178 1080 217
rect 1152 209 1231 217
rect 1152 182 1205 209
rect 1228 182 1231 209
rect 1152 178 1231 182
rect 628 151 673 178
rect -14 138 52 151
rect -14 98 1 138
rect 42 98 52 138
rect -14 80 52 98
rect 206 138 272 151
rect 206 98 220 138
rect 261 98 272 138
rect 206 80 272 98
rect 387 138 453 151
rect 387 98 402 138
rect 443 98 453 138
rect 387 80 453 98
rect 607 138 673 151
rect 607 98 621 138
rect 662 98 673 138
rect 607 80 673 98
rect 1548 116 1614 129
rect 1548 76 1563 116
rect 1604 76 1614 116
rect -14 49 52 62
rect -14 9 1 49
rect 42 9 52 49
rect -14 -9 52 9
rect 206 45 272 63
rect 387 49 453 62
rect 387 45 402 49
rect 206 43 402 45
rect 206 3 216 43
rect 257 9 402 43
rect 443 9 453 49
rect 257 3 453 9
rect 206 -3 453 3
rect 206 -8 272 -3
rect -310 -562 -278 -17
rect 213 -53 256 -8
rect 387 -9 453 -3
rect 607 43 673 63
rect 1548 58 1614 76
rect 1768 116 1834 129
rect 1768 76 1782 116
rect 1823 76 1834 116
rect 1768 58 1834 76
rect 607 3 617 43
rect 658 3 673 43
rect 607 -8 673 3
rect 1548 27 1614 40
rect 1548 -13 1563 27
rect 1604 -13 1614 27
rect 1548 -31 1614 -13
rect 1768 21 1834 41
rect 1768 -19 1778 21
rect 1819 -19 1834 21
rect 1768 -30 1834 -19
rect 87 -76 166 -60
rect 87 -114 99 -76
rect 146 -114 166 -76
rect -182 -127 -34 -119
rect -182 -197 -169 -127
rect -99 -197 -34 -127
rect -182 -208 -34 -197
rect 87 -160 166 -114
rect 87 -198 102 -160
rect 149 -198 166 -160
rect 87 -203 166 -198
rect 210 -171 256 -53
rect 494 -70 573 -52
rect 494 -108 512 -70
rect 559 -108 573 -70
rect 494 -149 573 -108
rect 274 -171 328 -169
rect 210 -199 328 -171
rect 494 -187 508 -149
rect 555 -187 573 -149
rect 494 -195 573 -187
rect 216 -205 328 -199
rect 274 -296 328 -205
rect 263 -309 329 -296
rect 263 -349 278 -309
rect 319 -349 329 -309
rect 263 -367 329 -349
rect -530 -967 -476 -953
rect -530 -998 -516 -967
rect -489 -989 -476 -967
rect -454 -981 -400 -967
rect -454 -989 -440 -981
rect -489 -998 -440 -989
rect -530 -1011 -440 -998
rect -530 -1027 -481 -1011
rect -454 -1012 -440 -1011
rect -413 -1012 -400 -981
rect -454 -1016 -400 -1012
rect -382 -978 -328 -964
rect -382 -1009 -368 -978
rect -341 -1009 -328 -978
rect -382 -1013 -328 -1009
rect -451 -1024 -400 -1016
rect -379 -1025 -328 -1013
rect -310 -1025 -279 -562
rect -254 -989 -215 -981
rect -254 -1020 -248 -989
rect -221 -1015 -215 -989
rect -221 -1016 -214 -1015
rect -221 -1020 -212 -1016
rect -254 -1025 -212 -1020
rect -379 -1050 -279 -1025
rect -256 -1048 -212 -1025
rect -373 -1053 -279 -1050
rect -369 -1054 -346 -1053
rect -249 -1084 -214 -1048
rect -248 -1140 -216 -1084
rect -270 -1153 -204 -1140
rect -270 -1193 -255 -1153
rect -214 -1193 -204 -1153
rect -270 -1211 -204 -1193
rect -282 -1829 -216 -1816
rect -282 -1869 -267 -1829
rect -226 -1869 -216 -1829
rect -282 -1887 -216 -1869
rect -62 -1829 4 -1816
rect -62 -1869 -48 -1829
rect -7 -1869 4 -1829
rect -62 -1887 4 -1869
rect 1548 -1886 1614 -1873
rect -282 -1918 -216 -1905
rect -282 -1958 -267 -1918
rect -226 -1958 -216 -1918
rect -282 -1976 -216 -1958
rect -62 -1924 4 -1904
rect -62 -1964 -52 -1924
rect -11 -1964 4 -1924
rect 1548 -1926 1563 -1886
rect 1604 -1926 1614 -1886
rect 1548 -1944 1614 -1926
rect 1768 -1886 1834 -1873
rect 1768 -1926 1782 -1886
rect 1823 -1926 1834 -1886
rect 1768 -1944 1834 -1926
rect -62 -1975 4 -1964
rect 252 -1969 318 -1956
rect -272 -2290 -230 -1976
rect 252 -2009 267 -1969
rect 308 -2009 318 -1969
rect 252 -2027 318 -2009
rect 472 -1969 538 -1956
rect 472 -2009 486 -1969
rect 527 -2009 538 -1969
rect 472 -2027 538 -2009
rect 1548 -1975 1614 -1962
rect 1548 -2015 1563 -1975
rect 1604 -2015 1614 -1975
rect 1548 -2033 1614 -2015
rect 1768 -1981 1834 -1961
rect 1768 -2021 1778 -1981
rect 1819 -2021 1834 -1981
rect 1768 -2032 1834 -2021
rect 252 -2058 318 -2045
rect 252 -2098 267 -2058
rect 308 -2098 318 -2058
rect 252 -2116 318 -2098
rect 472 -2064 538 -2044
rect 472 -2104 482 -2064
rect 523 -2104 538 -2064
rect 472 -2111 489 -2104
rect 507 -2111 538 -2104
rect 472 -2115 538 -2111
rect 342 -2267 1755 -2250
rect -176 -2268 1755 -2267
rect -176 -2283 1671 -2268
rect -176 -2290 367 -2283
rect -290 -2325 -161 -2290
rect -107 -2318 367 -2290
rect 421 -2301 1671 -2283
rect 1719 -2301 1755 -2268
rect 421 -2318 1755 -2301
rect -107 -2321 1755 -2318
rect -107 -2325 436 -2321
rect -290 -2337 436 -2325
rect -176 -2343 436 -2337
rect 1788 -2417 1811 -2032
rect 1701 -2456 1811 -2417
rect -135 -2459 1811 -2456
rect -135 -2498 -45 -2459
rect -23 -2471 1811 -2459
rect -23 -2498 492 -2471
rect 509 -2498 1811 -2471
rect -135 -2515 1811 -2498
<< viali >>
rect 217 1532 244 1552
rect 441 1536 468 1556
rect 219 1216 247 1238
rect 441 1216 469 1238
rect 1205 182 1228 209
rect 102 -198 149 -160
rect 508 -187 555 -149
rect -42 -1963 -23 -1941
rect 489 -2104 507 -2082
rect 489 -2111 507 -2104
rect -45 -2498 -23 -2459
rect 492 -2498 509 -2471
<< metal1 >>
rect 212 1552 254 1561
rect 212 1532 217 1552
rect 244 1532 254 1552
rect 212 1238 254 1532
rect 212 1216 219 1238
rect 247 1216 254 1238
rect 212 1209 254 1216
rect 434 1556 476 1561
rect 434 1536 441 1556
rect 468 1536 476 1556
rect 434 1238 476 1536
rect 434 1216 441 1238
rect 469 1216 476 1238
rect 434 1209 476 1216
rect 1198 209 1264 217
rect 1198 182 1205 209
rect 1228 182 1264 209
rect 1198 178 1264 182
rect 504 -149 561 -143
rect 98 -160 155 -152
rect 98 -198 102 -160
rect 149 -198 155 -160
rect 98 -217 155 -198
rect 504 -187 508 -149
rect 555 -180 561 -149
rect 555 -187 741 -180
rect 504 -208 741 -187
rect 507 -213 741 -208
rect -50 -1941 -15 -1930
rect -50 -1963 -42 -1941
rect -23 -1963 -15 -1941
rect -50 -2459 -15 -1963
rect -50 -2498 -45 -2459
rect -23 -2498 -15 -2459
rect -50 -2515 -15 -2498
rect 485 -2082 514 -2074
rect 485 -2111 489 -2082
rect 507 -2111 514 -2082
rect 485 -2471 514 -2111
rect 485 -2498 492 -2471
rect 509 -2498 514 -2471
rect 485 -2506 514 -2498
<< labels >>
rlabel metal1 1247 194 1247 194 1 out2
rlabel metal1 121 -211 121 -211 1 in1
rlabel locali 64 1534 64 1534 1 vdd
rlabel locali 815 -2490 815 -2490 1 vss
rlabel metal1 688 -197 688 -197 1 in2
rlabel locali -54 -173 -54 -173 1 vss
<< end >>
